module decoder (reg_in, decode_out);
input [4:0] reg_in;
output [31:0] decode_out;
 wire n_a, n_b, n_c, n_d, n_e;
 assign n_a = ~reg_in[4];
 assign n_b = ~reg_in[3];
 assign n_c = ~reg_in[2];
 assign n_d = ~reg_in[1];
 assign n_e = ~reg_in[0];
 and(decode_out[0], n_a, n_b, n_c, n_d, n_e);
 and(decode_out[1], n_a, n_b, n_c, n_d, reg_in[0]);
 and(decode_out[2], n_a, n_b, n_c, reg_in[1], n_e);
 and(decode_out[3], n_a, n_b, n_c, reg_in[1], reg_in[0]);
 and(decode_out[4], n_a, n_b, reg_in[2], n_d, n_e);
 and(decode_out[5], n_a, n_b, reg_in[2], n_d, reg_in[0]);
 and(decode_out[6], n_a, n_b, reg_in[2], reg_in[1], n_e);
 and(decode_out[7], n_a, n_b, reg_in[2], reg_in[1], reg_in[0]);
 and(decode_out[8], n_a, reg_in[3], n_c, n_d, n_e);
 and(decode_out[9], n_a, reg_in[3], n_c, n_d, reg_in[0]);
 and(decode_out[10], n_a, reg_in[3], n_c, reg_in[1], n_e);
 and(decode_out[11], n_a, reg_in[3], n_c,reg_in[1], reg_in[0]);
 and(decode_out[12], n_a, reg_in[3], reg_in[2], n_d, n_e);
 and(decode_out[13], n_a, reg_in[3], reg_in[2], n_d, reg_in[0]);
 and(decode_out[14], n_a, reg_in[3], reg_in[2], reg_in[1], n_e);
 and(decode_out[15], n_a, reg_in[3], reg_in[2], reg_in[1], reg_in[0]);
 and(decode_out[16], reg_in[4], n_b, n_c, n_d, n_e);
 and(decode_out[17], reg_in[4], n_b, n_c, n_d, reg_in[0]);
 and(decode_out[18], reg_in[4], n_b, n_c, reg_in[1], n_e);
 and(decode_out[19], reg_in[4], n_b, n_c, reg_in[1], reg_in[0]);
 and(decode_out[20], reg_in[4], n_b, reg_in[2], n_d, n_e);
 and(decode_out[21], reg_in[4], n_b, reg_in[2], n_d, reg_in[0]);
 and(decode_out[22], reg_in[4], n_b, reg_in[2], reg_in[1], n_e);
 and(decode_out[23], reg_in[4], n_b, reg_in[2], reg_in[1], reg_in[0]);
 and(decode_out[24], reg_in[4], reg_in[3], n_c, n_d, n_e);
 and(decode_out[25], reg_in[4], reg_in[3], n_c, n_d, reg_in[0]);
 and(decode_out[26], reg_in[4], reg_in[3], n_c, reg_in[1], n_e);
 and(decode_out[27], reg_in[4], reg_in[3], n_c, reg_in[1], reg_in[0]);
 and(decode_out[28], reg_in[4], reg_in[3], reg_in[2], n_d, n_e);
 and(decode_out[29], reg_in[4], reg_in[3], reg_in[2], n_d, reg_in[0]);
 and(decode_out[30], reg_in[4], reg_in[3], reg_in[2], reg_in[1], n_e);
 and(decode_out[31], reg_in[4], reg_in[3], reg_in[2], reg_in[1], reg_in[0]);

endmodule